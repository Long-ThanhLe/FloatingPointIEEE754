
module TAYLOR_EXP(
	in,
	out
);
input [31:0]in;
output [31:0]out;

// reg [32 -1 :0 ] num0375    = 32'b00111110110000000000000000000000;

// reg [32 -1 :0 ] num_ln0375 = 32'b1_01111110_11110110001011110100000;

// reg [32 -1 :0 ] num_ln2    = 32'b0_01111110_01100010111001000011000;

// wire [31:0] x_a_1;
// ADD X_A(.a(in[31:0]), .b(num0375[31:0]), .out(x_a_1[31:0]), .symbol(1'b1));

// wire [31:0] x_a_a_1;
// DIV X_A_A(.in1(x_a_1[31:0]), .in2(num0375[31:0]), .out(x_a_a_1[31:0]));
// DIV X_A_A(.in1(32'd0]), .in2(num0375[31:0]), .out(x_a_a_1[31:0]));

wire [31:0]  x_2, x_3, x_4, x_5, x_6;


MUL X_A_2(.in1(in[31:0]), .in2(in[31:0]), .out(x_2[31:0]));
MUL X_A_3(.in1(in[31:0]), .in2(x_2[31:0]), .out(x_3[31:0]));
MUL X_A_4(.in1(in[31:0]), .in2(x_3[31:0]), .out(x_4[31:0]));
MUL X_A_5(.in1(in[31:0]), .in2(x_4[31:0]), .out(x_5[31:0]));
MUL X_A_6(.in1(in[31:0]), .in2(x_5[31:0]), .out(x_6[31:0]));

wire [31:0] x__2, x__3, x__4, x__5, x__6;

DIV X_A_A__2(.in1(x_2[31:0]), .in2(32'b01000000000000000000000000000000), .out(x__2[31:0]));
DIV X_A_A__3(.in1(x_3[31:0]), .in2(32'b01000000110000000000000000000000), .out(x__3[31:0]));
DIV X_A_A__4(.in1(x_4[31:0]), .in2(32'b01000001110000000000000000000000), .out(x__4[31:0]));
DIV X_A_A__5(.in1(x_5[31:0]), .in2(32'b01000010111100000000000000000000), .out(x__5[31:0]));
DIV X_A_A__6(.in1(x_6[31:0]), .in2(32'b01000100001101000000000000000000), .out(x__6[31:0]));

wire [31:0] sum_1, sum_2,sum_3,sum_4,sum_5,sum_6;
ADD SUM_1 (.a(32'b00111111100000000000000000000000), .b(in[31:0]), .symbol(1'b0), .out(sum_1[31:0])  );
ADD SUM_2 (.a(sum_1[31:0]), .b(x__2[31:0]), .symbol(1'b0), .out(sum_2[31:0])  );
ADD SUM_3 (.a(sum_2[31:0]), .b(x__3[31:0]), .symbol(1'b0), .out(sum_3[31:0])  );
ADD SUM_4 (.a(sum_3[31:0]), .b(x__4[31:0]), .symbol(1'b0), .out(sum_4[31:0])  );
ADD SUM_5 (.a(sum_4[31:0]), .b(x__5[31:0]), .symbol(1'b0), .out(sum_5[31:0])  );
ADD SUM_6 (.a(sum_5[31:0]), .b(x__6[31:0]), .symbol(1'b0), .out(sum_6[31:0])  );

assign  out[31:0] = sum_6[31:0];

endmodule
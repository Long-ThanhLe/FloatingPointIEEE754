
module MUL_tb( );
	
reg [32-1:0]in1,in2;
wire[32-1:0]out;

MUL MUL_0(.in1(in1),.in2(in2),.out(out));
initial begin
	in1 = 32'b01000000000000000000000000000000;

	in2 = 32'b00111111100000000000000000000000;
	#10;

	in1 = 32'b01000000000000000000000000000000;

	in2 = 32'b01000000000000000000000000000000;
	#10;
	
	in1 = 32'b01000000101010000000000000000000;

	in2 = 32'b01000000000000000000000000000000;
	#10;
	in1 = 32'b10111111100000000000000000000000; //-1

	in2 = 32'b01000000000000000000000000000000;
	#10;
	in1 = 32'b01000000001000000000000000000000; //2.5

	in2 = 32'b01000000011000000000000000000000; //3.5
	#10;
	in1 = 32'b01000100111111000111001100110011; //2019.6
	
	in2 = 32'b11000000011000000000000000000000; //-3.5
	#10;

	in1 = 32'b01000100111111000111001100110011; //2019.6
	
	in2 = 32'b11111111100000000000000000000001;// NaN

	#10;
	in1 = 32'b0_00000000_00000000000000000000000; // 0
	
	in2 = 32'b0_00000000_00000000000000000000000; // 0

	#10;
	in1 = 32'b1_11111111_00000000000000000000000;// -INF
	
	in2 = 32'b0_11111111_00000000000000000000000;// +INF

	#10;
	in1 = 32'b0_11111111_00000000000000000000000;// +INF
	
	in2 = 32'b0_00000000_00000000000000000000000;// 0

	#10;
	in1 = 32'b1_11111111_00000000000000000000000;// -INF
	
	in2 = 32'b1_11111111_00000000000000000000000;// -INF

	#10;
	in1 = 32'b0_11111111_00000000000000000000000;// +INF
	
	in2 = 32'b1_11111111_00000000000000000000000;// -INF



end
	
endmodule 
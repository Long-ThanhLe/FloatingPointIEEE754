module ADD(
    a,
    b,
    symbol,
    out
);

endmodule

module MUL_tb( );
	
reg [32-1:0]in1,in2;
wire[32-1:0]out;

MUL MUL_0(.in1(in1),.in2(in2),.out(out));
initial begin
	#10;
	in1 = 32'b01000000000000000000000000000000;

	in2 = 32'b00111111100000000000000000000000;
	#10;

	in1 = 32'b01000000000000000000000000000000;

	in2 = 32'b01000000000000000000000000000000;
	#10;
	
	in1 = 32'b01000000101010000000000000000000;

	in2 = 32'b01000000000000000000000000000000;
	#10;
	
end
	
endmodule 
module ADD_tb();

parameter DATA_WIDTH = 32;

reg   [DATA_WIDTH - 1:  0]  a, b;
reg   symbol;
wire  [DATA_WIDTH - 1: 0] out;

ADD     ADD_TB(.a(a),   .b(b),  .symbol(symbol), .out(out));

initial
begin
  a = 32'b01000000101000000000000000000000;
  b = 32'b01000000111000000000000000000000;
  symbol = 0;
  #10;
  a = 32'b01000000101000000000000000000000;
  b = 32'b01000000111000000000000000000000;
  symbol = 1;
  #10;
  a = 32'b00000000000000000000000000000000; //-15.6
  b = 32'b01000000011011001100110011001101; // 3.7
  symbol = 0;
  #10;
  a = 32'b11000001011110011001100110011010; //-15.6
  b = 32'b01000000011011001100110011001101; // 3.7
  symbol = 1;
  #10;
  a = 32'b11000001011110011001100110011010; // 15.6
  b = 32'b11000000011011001100110011001101; // 3.7
  symbol = 0;
  #10;
  #10;
  a = 32'b0_01111101_10000000000000000000000; // 0.375
  b = 32'b0_01111101_10000000000000000000000; // 0.375
  symbol = 1'b1;
end


endmodule
module CONVERTER_BI_2_DEC_tb();

reg [31:0]in;
wire [127:0]out_floor, out_frac;
wire out_sign;

COVERT_BI_2_DEC CONV(.in(in), .out_floor(out_floor), .out_frac(out_frac), .out_sign(out_sign));

initial begin

	#10;
	in = 32'b01000000000000000000000000000000;//2
	#10;
	in = 32'b01000000010000000000000000000000;//3
	#10;
	in = 32'b01000000011001100110011001100110;//3.6
	#10;
	in = 32'b01000010011000000000000000110100;//56.0002
	#10;
	in = 32'b01000010110010000110011001100110;//100.2
	#10;
	in = 32'b00111001010100011011011100010111;//0.0002
	#10;
	in = 32'b00111100101000111101011100001010;//0.02
	#10;
	in = 32'b00111110010011001100110011001101;//0.2
	#10;
	in = 32'b01000000010000000101000111101100;//3.005
	#10;
	in = 32'b01000010011000000000000000110100;//56.0002
end
endmodule

